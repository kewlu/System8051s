----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Thu May 11 13:22:17 2017
-- Parameters for CoreTimer
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant FAMILY : integer := 16;
    constant INTACTIVEH : integer := 1;
    constant WIDTH : integer := 32;
end coreparameters;
